// alu.v
// RV32I ALU supporting arithmetic, logic, and shift operations.
`timescale 1ns/1ps

module alu (
    input      [31:0] op_a,
    input      [31:0] op_b,
    input      [3:0]  alu_ctrl,
    output reg [31:0] result,
    output            zero
);
    localparam ALU_ADD  = 4'b0000;
    localparam ALU_SUB  = 4'b0001;
    localparam ALU_AND  = 4'b0010;
    localparam ALU_OR   = 4'b0011;
    localparam ALU_XOR  = 4'b0100;
    localparam ALU_SLT  = 4'b0101;
    localparam ALU_SLTU = 4'b0110;
    localparam ALU_SLL  = 4'b0111;
    localparam ALU_SRL  = 4'b1000;
    localparam ALU_SRA  = 4'b1001;

    always @(*) begin
        case (alu_ctrl)
            ALU_ADD:  result = op_a + op_b;
            ALU_SUB:  result = op_a - op_b;
            ALU_AND:  result = op_a & op_b;
            ALU_OR:   result = op_a | op_b;
            ALU_XOR:  result = op_a ^ op_b;
            ALU_SLT:  result = ($signed(op_a) < $signed(op_b)) ? 32'h1 : 32'h0;
            ALU_SLTU: result = (op_a < op_b) ? 32'h1 : 32'h0;
            ALU_SLL:  result = op_a << op_b[4:0];
            ALU_SRL:  result = op_a >> op_b[4:0];
            ALU_SRA:  result = $signed(op_a) >>> op_b[4:0];
            default:  result = 32'h0;
        endcase
    end

    assign zero = (result == 32'h0);
endmodule
